`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:26:13 12/15/2022 
// Design Name: 
// Module Name:    ALU_Main 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALU_Main(
    input [15:0] data_in_1,
    input [15:0] data_in_2,
    input [1:0] alu_op,
    output [15:0] data_out,
    output z_flag,
    output a_grt_b,
    output b_grt_a
    );
	 
	 
	 


endmodule
